* LM311 VOLTAGE COMPARATOR "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS VERSION 4.03 ON 03/07/90 AT 08:15
* REV (N/A)
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OPEN COLLECTOR OUTPUT
*                | | | | | OUTPUT GROUND
*                | | | | | |
.SUBCKT LM311    1 2 3 4 5 6
*
  F1    9  3 V1 1
  IEE   3  7 DC 100.0E-6
  VI1  21  1 DC .45
  VI2  22  2 DC .45
  Q1    9 21  7 QIN
  Q2    8 22  7 QIN
  Q3    9  8  4 QMO
  Q4    8  8  4 QMI
.MODEL QIN PNP(IS=800.0E-18 BF=500)
.MODEL QMI NPN(IS=800.0E-18 BF=1002)
.MODEL QMO NPN(IS=800.0E-18 BF=1000 CJC=1E-15 TR=102.5E-9)
  E1   10  6  9  4  1
  V1   10 11 DC 0
  Q5    5 11  6 QOC
.MODEL QOC NPN(IS=800.0E-18 BF=103.5E3 CJC=1E-15 TF=11.60E-12 TR=48.19E-9)
  DP    4  3 DX
  RP    3  4 6.667E3
.MODEL DX  D(IS=800.0E-18)
.ENDS
